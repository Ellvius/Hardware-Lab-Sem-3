module BCD_counter();

endmodule

