module Custom_register();

endmodule
