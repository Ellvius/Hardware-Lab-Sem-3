module BCD_counter_tb;

endmodule

