
module Sequence_detector();
endmodule
