module Vending_machine();
endmodule
