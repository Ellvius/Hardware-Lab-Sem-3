module Vending_machine_tb;
endmodule
