module Updown_synchronous_counter();

endmodule
