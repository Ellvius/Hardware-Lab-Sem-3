module Updown_synchronous_counter_tb;

endmodule
