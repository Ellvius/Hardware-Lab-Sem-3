module SIPO();

endmodule
