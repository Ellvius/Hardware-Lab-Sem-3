module SIPO_tb;

endmodule
