module Custom_register_tb;

endmodule
