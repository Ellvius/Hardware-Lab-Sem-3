module Sequence_detector_tb;
endmodule
